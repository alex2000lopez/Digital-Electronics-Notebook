entity NAME_ENTITY is
    port(NAME_OF_PORT_1:  DIRECTION  DATA_TYPE;
                        . . .
         );
  end NAME_ENTITY;