architecture ARCH of NAME_ENTITY is
    --begin
    --  process(sensitivity list)
      begin
        concurrent/sequential instructions
    end ARCH;